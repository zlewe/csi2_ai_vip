interface csi2_if (input bit clk); // 'clk' is a general system clock or reference clock

    // D-PHY related signals (simplified for driver interaction)
    // The actual differential pairs (p/n) and tristate buffers would be instantiated
    // at a lower level or within the interface's internal logic, mapping these
    // abstract byte/bit signals to physical wires.

    // High-speed Lane Clock Input: This clock is typically generated by the PHY
    // or a dedicated clock generator and used by the driver for synchronization.
    logic hs_lane_clk_i;

    // High-speed Data Lanes (up to 4 lanes):
    // 'hs_data_out' represents the byte data driven on each lane.
    // 'hs_data_oe' controls the output enable for each lane's high-speed data drivers.
    logic [7:0] hs_data_out[3:0]; // Output byte data for up to 4 lanes
    logic       hs_data_oe[3:0];  // Output enable for high-speed data lanes (1 per lane)

    // High-speed Clock Lane:
    // 'hs_clk_out' represents the high-speed clock signal (e.g., continuous clock in D-PHY).
    // 'hs_clk_oe' controls the output enable for the high-speed clock driver.
    logic hs_clk_out;             // Output clock signal
    logic hs_clk_oe;              // Output enable for high-speed clock lane

    // Low-power Mode Control Signals:
    // These signals control the transition between high-speed and low-power modes.
    logic lp_mode_en[3:0];        // Enable low-power mode per data lane (1: LP, 0: HS)
    logic lp_mode_clk_en;         // Enable low-power mode for clock lane (1: LP, 0: HS)

    // Low-power Data/Clock (used for control/escape mode commands)
    logic [7:0] lp_data_out[3:0]; // Output data in low-power mode (e.g., for escape sequences)
    logic       lp_data_oe[3:0];  // Output enable for low-power data lanes
    logic lp_clk_out;             // Output clock in low-power mode
    logic lp_clk_oe;              // Output enable for low-power clock lane

    // Reset signal (driven by driver)
    logic reset_n_out;            // Active low reset signal
    logic reset_n_oe;             // Output enable for reset signal

    // Modport for the Driver
    // Defines the signals that the `csi2_driver` can control or observe.
    modport driver_mp (
        // Outputs controlled by the driver
        output hs_data_out,       // Array of 4 bytes
        output hs_data_oe,        // Array of 4 bits
        output hs_clk_out,
        output hs_clk_oe,
        output lp_mode_en,        // Array of 4 bits
        output lp_mode_clk_en,
        output lp_data_out,       // Array of 4 bytes
        output lp_data_oe,        // Array of 4 bits
        output lp_clk_out,
        output lp_clk_oe,
        output reset_n_out,
        output reset_n_oe,
        // Inputs observed by the driver (e.g., for timing synchronization)
        input hs_lane_clk_i
    );

    // Modport for the Monitor (or other components observing the interface)
    // Defines the signals that a `csi2_monitor` would observe.
    modport monitor_mp (
        input hs_data_out,
        input hs_data_oe,
        input hs_clk_out,
        input hs_clk_oe,
        input lp_mode_en,
        input lp_mode_clk_en,
        input lp_data_out,
        input lp_data_oe,
        input lp_clk_out,
        input lp_clk_oe,
        input reset_n_out,
        input reset_n_oe,
        input hs_lane_clk_i
    );

endinterface
